/*-----------------------------------------------------------------------
				shift rows transformation
-----------------------------------------------------------------------*/
module Shift_Rows_Enc
	(
	input  [127:0] i_Din, // Data input to be transformed
	output [127:0] o_Dout
	);
assign o_Dout[007:000] = i_Din[039:032];// As the high data are put into the situation of 0//
assign o_Dout[015:008] = i_Din[079:072]; // So o_Dout[127:120] represent for 0 byte which is in the poly.//
assign o_Dout[023:016] = i_Din[119:112];
assign o_Dout[031:024] = i_Din[031:024];
assign o_Dout[039:032] = i_Din[071:064];
assign o_Dout[047:040] = i_Din[111:104];
assign o_Dout[055:048] = i_Din[023:016];
assign o_Dout[063:056] = i_Din[063:056];
assign o_Dout[071:064] = i_Din[103:096];
assign o_Dout[079:072] = i_Din[015:008];
assign o_Dout[087:080] = i_Din[055:048];
assign o_Dout[095:088] = i_Din[095:088];
assign o_Dout[103:096] = i_Din[007:000];
assign o_Dout[111:104] = i_Din[047:040];
assign o_Dout[119:112] = i_Din[087:080];
assign o_Dout[127:120] = i_Din[127:120];
endmodule